
library ieee;
use ieee.std_logic_1164.all;

library surf;
use surf.StdRtlPkg.all;
use surf.AxiLitePkg.all;

-------------------------------------------------------------------------------
-- File       : AppPkg.vhd
-- Company    : SLAC National Accelerator Laboratory
-------------------------------------------------------------------------------
-- Description: Application's Package File
-------------------------------------------------------------------------------
-- This file is part of 'EPIX HR Firmware'.
-- It is subject to the license terms in the LICENSE.txt file found in the 
-- top-level directory of this distribution and at: 
--    https://confluence.slac.stanford.edu/display/ppareg/LICENSE.html. 
-- No part of 'EPIX HR Firmware', including this file, 
-- may be copied, modified, propagated, or distributed except according to 
-- the terms contained in the LICENSE.txt file.
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

library surf;
use surf.StdRtlPkg.all;
use surf.AxiLitePkg.all;

package AppPkg is

   constant XIL_DEVICE_C                    : string  := "ULTRASCALE_PLUS";
   constant NUMBER_OF_ASICS_C               : natural := 4;   
   constant NUMBER_OF_LANES_C               : natural := 1;

   constant NUM_AXIL_MASTERS_C              : natural := 1;
   constant NUM_AXIL_SLAVES_C               : natural := 1;

   constant PLLREGS_AXI_INDEX_C             : natural := 0;
   constant PLLREGS_AXI_BASE_ADDR_C         : slv(31 downto 0) := X"80000000";--0 
   
   -- constant XBAR_CONFIG_C : AxiLiteCrossbarMasterConfigArray(NUM_AXIL_MASTERS_C-1 downto 0) := (
   --    PLLREGS_AXI_INDEX_C       => (
   --       baseAddr             => PLLREGS_AXI_BASE_ADDR_C,
   --       addrBits             => 24,
   --       connectivity         => x"FFFF"));


   

end package AppPkg;

package body AppPkg is

end package body AppPkg;
